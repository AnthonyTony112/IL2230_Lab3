library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.fixed_pkg.all;

entity nonlinear is
	generic (int_bit: integer :=3; float_bit: integer := 5);
	port (
		output: IN sfixed (int_bit-1 downto -float_bit);
		Reluout: Out sfixed (int_bit-1 downto -float_bit)
		--sigout: Out std_logic_vector (int_bit+float_bit-1 downto 0)
	);
end nonlinear;

architecture behave of nonlinear is
    subtype Data is std_logic_vector(int_bit+float_bit-1 downto 0);
    signal input : std_logic_vector (int_bit+float_bit-1 downto 0):=(others=>'0');
--    type LUTArray is array(0 to 255) of Data;
--    signal index : std_logic_vector(7 downto 0):="00000000";
--	signal inputpre: sfixed(int_bit-1 downto -float_bit):=(0=>'1',others=>'0');
--	signal indexin: integer:=0;
    constant one: sfixed(int_bit-1 downto -float_bit):=(0=>'1',others=>'0');
    constant clamp: std_logic_vector((int_bit+float_bit-1) downto 0) := ((int_bit+float_bit-1) => '0', others => '1');
    constant zeroR: sfixed (int_bit-1 downto -float_bit):=(others=>'0');
--    constant LUTSigmoid :LUTArray:=(
--		x"00",
--		x"00",
--		x"00",
--		x"00",
--		x"00",
--		x"00",
--		x"00",
--		x"00",
--		x"00",
--		x"00",
--		x"00",
--		x"00",
--		x"00",
--		x"00",
--		x"00",
--		x"00",
--		x"00",
--		x"00",
--		x"00",
--		x"01",
--		x"01",
--		x"01",
--		x"01",
--		x"01",
--		x"01",
--		x"01",
--		x"01",
--		x"01",
--		x"01",
--		x"01",
--		x"01",
--		x"01",
--		x"01",
--		x"01",
--		x"01",
--		x"01",
--		x"01",
--		x"01",
--		x"01",
--		x"01",
--		x"01",
--		x"01",
--		x"02",
--		x"02",
--		x"02",
--		x"02",
--		x"02",
--		x"02",
--		x"02",
--		x"02",
--		x"02",
--		x"02",
--		x"02",
--		x"02",
--		x"02",
--		x"02",
--		x"03",
--		x"03",
--		x"03",
--		x"03",
--		x"03",
--		x"03",
--		x"03",
--		x"03",
--		x"03",
--		x"03",
--		x"04",
--		x"04",
--		x"04",
--		x"04",
--		x"04",
--		x"04",
--		x"04",
--		x"04",
--		x"05",
--		x"05",
--		x"05",
--		x"05",
--		x"05",
--		x"05",
--		x"05",
--		x"06",
--		x"06",
--		x"06",
--		x"06",
--		x"06",
--		x"06",
--		x"07",
--		x"07",
--		x"07",
--		x"07",
--		x"07",
--		x"07",
--		x"08",
--		x"08",
--		x"08",
--		x"08",
--		x"08",
--		x"09",
--		x"09",
--		x"09",
--		x"09",
--		x"09",
--		x"0A",
--		x"0A",
--		x"0A",
--		x"0A",
--		x"0B",
--		x"0B",
--		x"0B",
--		x"0B",
--		x"0B",
--		x"0C",
--		x"0C",
--		x"0C",
--		x"0C",
--		x"0D",
--		x"0D",
--		x"0D",
--		x"0D",
--		x"0E",
--		x"0E",
--		x"0E",
--		x"0E",
--		x"0F",
--		x"0F",
--		x"0F",
--		x"0F",
--		x"10",
--		x"10",
--		x"10",
--		x"10",
--		x"11",
--		x"11",
--		x"11",
--		x"11",
--		x"12",
--		x"12",
--		x"12",
--		x"12",
--		x"13",
--		x"13",
--		x"13",
--		x"13",
--		x"14",
--		x"14",
--		x"14",
--		x"14",
--		x"14",
--		x"15",
--		x"15",
--		x"15",
--		x"15",
--		x"16",
--		x"16",
--		x"16",
--		x"16",
--		x"16",
--		x"17",
--		x"17",
--		x"17",
--		x"17",
--		x"17",
--		x"18",
--		x"18",
--		x"18",
--		x"18",
--		x"18",
--		x"18",
--		x"19",
--		x"19",
--		x"19",
--		x"19",
--		x"19",
--		x"19",
--		x"1A",
--		x"1A",
--		x"1A",
--		x"1A",
--		x"1A",
--		x"1A",
--		x"1A",
--		x"1B",
--		x"1B",
--		x"1B",
--		x"1B",
--		x"1B",
--		x"1B",
--		x"1B",
--		x"1B",
--		x"1C",
--		x"1C",
--		x"1C",
--		x"1C",
--		x"1C",
--		x"1C",
--		x"1C",
--		x"1C",
--		x"1C",
--		x"1C",
--		x"1D",
--		x"1D",
--		x"1D",
--		x"1D",
--		x"1D",
--		x"1D",
--		x"1D",
--		x"1D",
--		x"1D",
--		x"1D",
--		x"1D",
--		x"1D",
--		x"1D",
--		x"1D",
--		x"1E",
--		x"1E",
--		x"1E",
--		x"1E",
--		x"1E",
--		x"1E",
--		x"1E",
--		x"1E",
--		x"1E",
--		x"1E",
--		x"1E",
--		x"1E",
--		x"1E",
--		x"1E",
--		x"1E",
--		x"1E",
--		x"1E",
--		x"1E",
--		x"1E",
--		x"1E",
--		x"1E",
--		x"1E",
--		x"1E",
--		x"1F",
--		x"1F",
--		x"1F",
--		x"1F",
--		x"1F",
--		x"1F",
--		x"1F",
--		x"1F",
--		x"1F",
--		x"1F",
--		x"1F",
--		x"1F",
--		x"1F",
--		x"1F",
--		x"1F",
--		x"1F",
--		x"1F",
--		x"1F",
--		x"1F"		
--	--others=>"00000000"
--);
begin
	reluout <=zeroR when output<=zeroR else output;
--	inputpre<=output;
--	input<=to_slv(inputpre);
--	process(input)
--	  variable LUT_index : integer;
--		begin
--			if(int_bit>=4) then
--		 		sigout<=(others=>'0');
--		 	else
--				--input<=to_slv(output);
--				--input<="01101111";
--		 		if(signed(input) <= -signed(clamp)-1) then sigout <= LUTSigmoid(0);
--		 		elsif(signed(input) >= signed(clamp)) then sigout <= LUTSigmoid(2**6-1);
--		 		else 
--				 	--index<=std_logic_vector(signed(input)+signed(clamp));
--					--LUT_index := to_integer(unsigned(index));
--					LUT_index := to_integer(signed(input));
--					indexin<=to_integer(signed(input)); 
--					sigout <= LUTSigmoid(128+LUT_index);
--		 		end if;
--			end if;
--		 		
--       end process;
end behave; 


