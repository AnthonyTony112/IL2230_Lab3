library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.fixed_pkg.all;

entity nonlinear is
	generic (int_bit: integer :=6; float_bit: integer := 10);
	port (
		output: IN sfixed (int_bit-1 downto -float_bit);
		Reluout: Out sfixed (int_bit-1 downto -float_bit);
		sigout: Out sfixed (int_bit-1 downto -float_bit)
	);
end nonlinear;

architecture behave of nonlinear is
	subtype DataLUT is sfixed (2 downto -5);
    signal input : std_logic_vector (int_bit+float_bit-1 downto 0):=(others=>'0');
    type LUTArray is array(0 to 255) of DataLUT;
    signal index : std_logic_vector(7 downto 0):="00000000";
	signal inputpre: sfixed(int_bit-1 downto -float_bit):=(0=>'1',others=>'0');
	signal indexin: integer:=0;
    constant one: sfixed(int_bit-1 downto -float_bit):=(0=>'1',others=>'0');
    constant clamp: std_logic_vector((int_bit+float_bit-1) downto 0) := ((int_bit+float_bit-1) => '0', others => '1');
    constant zeroR: sfixed (int_bit-1 downto -float_bit):=(others=>'0');
    constant LUTSigmoid :LUTArray:=(
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000001",
		"00000001",
		"00000001",
		"00000001",
		"00000001",
		"00000001",
		"00000001",
		"00000001",
		"00000001",
		"00000001",
		"00000001",
		"00000001",
		"00000001",
		"00000001",
		"00000001",
		"00000001",
		"00000001",
		"00000001",
		"00000001",
		"00000001",
		"00000001",
		"00000001",
		"00000001",
		"00000010",
		"00000010",
		"00000010",
		"00000010",
		"00000010",
		"00000010",
		"00000010",
		"00000010",
		"00000010",
		"00000010",
		"00000010",
		"00000010",
		"00000010",
		"00000010",
		"00000011",
		"00000011",
		"00000011",
		"00000011",
		"00000011",
		"00000011",
		"00000011",
		"00000011",
		"00000011",
		"00000011",
		"00000100",
		"00000100",
		"00000100",
		"00000100",
		"00000100",
		"00000100",
		"00000100",
		"00000100",
		"00000101",
		"00000101",
		"00000101",
		"00000101",
		"00000101",
		"00000101",
		"00000101",
		"00000110",
		"00000110",
		"00000110",
		"00000110",
		"00000110",
		"00000110",
		"00000111",
		"00000111",
		"00000111",
		"00000111",
		"00000111",
		"00000111",
		"00001000",
		"00001000",
		"00001000",
		"00001000",
		"00001000",
		"00001001",
		"00001001",
		"00001001",
		"00001001",
		"00001001",
		"00001010",
		"00001010",
		"00001010",
		"00001010",
		"00001011",
		"00001011",
		"00001011",
		"00001011",
		"00001011",
		"00001100",
		"00001100",
		"00001100",
		"00001100",
		"00001101",
		"00001101",
		"00001101",
		"00001101",
		"00001110",
		"00001110",
		"00001110",
		"00001110",
		"00001111",
		"00001111",
		"00001111",
		"00001111",
		"00010000",
		"00010000",
		"00010000",
		"00010000",
		"00010001",
		"00010001",
		"00010001",
		"00010001",
		"00010010",
		"00010010",
		"00010010",
		"00010010",
		"00010011",
		"00010011",
		"00010011",
		"00010011",
		"00010100",
		"00010100",
		"00010100",
		"00010100",
		"00010100",
		"00010101",
		"00010101",
		"00010101",
		"00010101",
		"00010110",
		"00010110",
		"00010110",
		"00010110",
		"00010110",
		"00010111",
		"00010111",
		"00010111",
		"00010111",
		"00010111",
		"00011000",
		"00011000",
		"00011000",
		"00011000",
		"00011000",
		"00011000",
		"00011001",
		"00011001",
		"00011001",
		"00011001",
		"00011001",
		"00011001",
		"00011010",
		"00011010",
		"00011010",
		"00011010",
		"00011010",
		"00011010",
		"00011010",
		"00011011",
		"00011011",
		"00011011",
		"00011011",
		"00011011",
		"00011011",
		"00011011",
		"00011011",
		"00011100",
		"00011100",
		"00011100",
		"00011100",
		"00011100",
		"00011100",
		"00011100",
		"00011100",
		"00011100",
		"00011100",
		"00011101",
		"00011101",
		"00011101",
		"00011101",
		"00011101",
		"00011101",
		"00011101",
		"00011101",
		"00011101",
		"00011101",
		"00011101",
		"00011101",
		"00011101",
		"00011101",
		"00011110",
		"00011110",
		"00011110",
		"00011110",
		"00011110",
		"00011110",
		"00011110",
		"00011110",
		"00011110",
		"00011110",
		"00011110",
		"00011110",
		"00011110",
		"00011110",
		"00011110",
		"00011110",
		"00011110",
		"00011110",
		"00011110",
		"00011110",
		"00011110",
		"00011110",
		"00011110",
		"00011111",
		"00011111",
		"00011111",
		"00011111",
		"00011111",
		"00011111",
		"00011111",
		"00011111",
		"00011111",
		"00011111",
		"00011111",
		"00011111",
		"00011111",
		"00011111",
		"00011111",
		"00011111",
		"00011111",
		"00011111",
		"00011111"
	--others=>"00000000"
);
begin
	reluout <=zeroR when output<=zeroR else output;
	inputpre<=output;
	input<=to_slv(inputpre);
	process(input)
	  variable LUT_index : integer;
		begin
			if(int_bit>=4) then
		 		sigout<=(others=>'0');
		 	else
				--input<=to_slv(output);
				--input<="01101111";
		 		if(signed(input) <= -signed(clamp)-1) then sigout <= LUTSigmoid(0);
		 		elsif(signed(input) >= signed(clamp)) then sigout <= LUTSigmoid(2**6-1);
		 		else 
				 	--index<=std_logic_vector(signed(input)+signed(clamp));
					--LUT_index := to_integer(unsigned(index));
					LUT_index := to_integer(signed(input));
					indexin<=to_integer(signed(input)); 
					sigout <= LUTSigmoid(128+LUT_index);
		 		end if;
			end if;
		 		
       end process;
end behave; 


