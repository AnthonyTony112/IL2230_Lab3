library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.fixed_pkg.all;
USE work.all  ; 
USE work.CoeffPak.all  ; 
use IEEE.math_real.ceil;
use IEEE.math_real.log2;

entity ROM is
generic (
		N: integer:=3;
		M: integer:=3;
		int_bit: integer:=3;
		float_bit: integer:=5	
	);

port(addr: in std_logic_vector (7 downto 0);
     clk: in std_logic; 
     W: out DataArray2D);
end ROM;

architecture behave of ROM is
  
--signal W1D: DataArray
--type WeightArray is array(0 to 15) of sfixed (int_bit-1 downto -float_bit);
--type WeightArray2D is array (0 to 15) of WeightArray;
--type WeightArray3D is array (0 to 15) of WeightArray2D;
Constant Weight: DataArray3D:=

(

( 
  ("00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001"),
   
   ("00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010"),

   ("00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100"),

  ("00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001"),
   
   ("00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010"),

   ("00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100"),
    

  ("00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001"),
   
   ("00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010"),

   ("00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100"),
    
    ("00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001"),
   
   ("00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010"),

   ("00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100"),

  ("00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001"),
   
   ("00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010"),

   ("00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100"),
    

  ("00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001")
) , --layer1



( 
  ("00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001"),
   
   ("00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010"),

   ("00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100"),

  ("00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001"),
   
   ("00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010"),

   ("00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100"),
    

  ("00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001"),
   
   ("00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010"),

   ("00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100"),
    
    ("00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001"),
   
   ("00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010"),

   ("00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100"),

  ("00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001"),
   
   ("00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010"),

   ("00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100"),
    

  ("00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001")
) , --layer0

( 
  ("00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001"),
   
   ("00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010"),

   ("00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100"),

  ("00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001"),
   
   ("00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010"),

   ("00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100"),
    

  ("00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001"),
   
   ("00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010"),

   ("00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100"),
    
    ("00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001"),
   
   ("00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010"),

   ("00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100"),

  ("00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001"),
   
   ("00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010"),

   ("00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100"),
    

  ("00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001",
   "00000001")
) , --layer2



others=>(others=>(others=>(others=>'0')))
);
     
begin
  W<=Weight(to_integer(unsigned(addr)));

end behave;